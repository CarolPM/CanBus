module teste
reg test = 5'b01;
initial
    begin
		$display("%b", test);
	 end
   
endmodule